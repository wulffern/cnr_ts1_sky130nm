*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/CNR_TS1_lpe.spi
#else
.include ../../../work/lpe/SUN_PLL_ROSC_lpe.spi
.include ../../../work/xsch/CNR_TS1.spice

#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-4

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0
VDD  VDD_1V8  VSS  pwl 0 0 10n {AVDD}
VPWR  PWRUP_1V8  VSS  pwl 0 0 39n 0 40n {AVDD}

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
.include ../xdut.spi

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#endif
.save i(vdd)
.save v(do_1v8)
.save v(XDUT.VB_FVF) v(XDUT.VDD_ROSC) v(XDUT.VD)
.save v(PWRUP_1V8)
.save v(RST_N_1V8)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 10n 1u 0



foreach vtemp -40 -20 0 20 40 80 125

  option temp=$vtemp
  tran 1n 200n

  set fend = .raw
  write {cicname}_$vtemp$fend
end



quit


.endc

.end
