* NGSPICE file created from SUN_PLL_ROSC.ext - technology: sky130B

* Replacing the lpe port list (../tech/scripts/fixlpe)
.subckt SUN_PLL_ROSC AVDD CK VDD_ROSC PWRUP_1V8 AVSS
*.subckt SUN_PLL_ROSC CK PWRUP_1V8 VDD_ROSC AVDD AVSS
X0 CK xa3.YN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X1 CK xa3.YN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X2 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=11.6964 ps=62.7 w=1.08 l=0.18
X3 AVDD AVDD AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=3.6936 ps=19.8 w=1.08 l=0.18
X4 xa3.xc1b.S xa3.YN AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X5 xb2_3.Y xb2_2.Y VDD_ROSC AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X6 xb2_4.Y xb2_3.Y VDD_ROSC AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X7 xb2_3.Y xb2_2.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X8 xb2_4.Y xb2_3.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X9 xa3.Y xa3.AN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X10 xa3.Y xa3.YN xa3.xc1b.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X11 xa3.Y xa3.AN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X12 VDD_ROSC xb1.B xb2_0.A AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X13 xb2_0.A PWRUP_1V8 VDD_ROSC AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X14 xb2_0.A xb1.B xb1.MN1.S AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X15 xa3.YN xa3.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X16 xa3.xc2b.S xa3.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X17 xa3.AN xa3.A VDD_ROSC AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X18 xa3.A xb2_4.Y VDD_ROSC AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X19 xb2_0.Y xb2_0.A VDD_ROSC AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X20 xa3.AN xa3.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X21 xa3.A xb2_4.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X22 xb2_0.Y xb2_0.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X23 xa3.YN xa3.A AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X24 xa3.YN xa3.Y xa3.xc2b.S AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X25 xa4.Y xa3.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X26 xa4.Y xa3.Y AVDD AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X27 xb1.MN1.S PWRUP_1V8 AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X28 xb2_1.Y xb2_0.Y VDD_ROSC AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X29 xb3.MP1.G xb3.MP1.G xb3.MP1.G AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=1.2312 ps=6.6 w=1.08 l=0.18
X30 xb1.B xa3.AN VDD_ROSC AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X31 xb2_2.Y xb2_1.Y VDD_ROSC AVDD sky130_fd_pr__pfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X32 xb2_1.Y xb2_0.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X33 AVSS AVSS AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0 ps=0 w=1.08 l=0.18
X34 xb1.B xa3.AN AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
X35 xb2_2.Y xb2_1.Y AVSS AVSS sky130_fd_pr__nfet_01v8 ad=0.6156 pd=3.3 as=0.6156 ps=3.3 w=1.08 l=0.18
C0 a_2244_1454# AVDD 0.382164f
C1 xb2_4.Y xb2_3.Y 0.196604f
C2 xb2_0.A VDD_ROSC 0.226376f
C3 xb2_4.Y a_4764_3214# 0.126366f
C4 xb2_0.A AVDD 0.636038f
C5 a_3612_1806# AVDD 0.352245f
C6 a_2244_1806# AVDD 0.363881f
C7 xb2_0.Y VDD_ROSC 0.174397f
C8 xb2_0.Y AVDD 0.549611f
C9 xa3.xc2b.S AVDD 0.158852f
C10 xa3.A xb2_4.Y 0.227933f
C11 xa3.A a_4764_3566# 0.133585f
C12 a_3612_2158# AVDD 0.352242f
C13 a_2244_2158# AVDD 0.383825f
C14 xb2_0.A xb1.MN1.S 0.106429f
C15 xb2_1.Y VDD_ROSC 0.174326f
C16 xb2_1.Y AVDD 0.542798f
C17 xb2_0.A a_4764_1454# 0.126526f
C18 xa3.Y AVDD 1.88477f
C19 xa3.AN xa3.A 1.04758f
C20 xa4.Y AVDD 0.226929f
C21 xa3.AN a_4764_3918# 0.133315f
C22 a_3612_2510# AVDD 0.352239f
C23 a_2244_2510# AVDD 0.388264f
C24 xb1.B xa3.AN 0.19372f
C25 xb2_2.Y VDD_ROSC 0.174326f
C26 xb2_2.Y AVDD 0.542798f
C27 xa3.YN AVDD 1.81675f
C28 xb2_0.Y xb2_0.A 0.18371f
C29 a_3612_2862# AVDD 0.352239f
C30 xb2_0.Y a_4764_1806# 0.126366f
C31 a_2244_2862# AVDD 0.468641f
C32 xb2_3.Y VDD_ROSC 0.174326f
C33 xb2_3.Y AVDD 0.545348f
C34 a_3612_3214# AVDD 0.351928f
C35 xa3.Y a_2244_1454# 0.113253f
C36 a_2244_3214# AVDD 0.439118f
C37 xa3.YN a_2244_1102# 0.164472f
C38 xb2_4.Y VDD_ROSC 0.173007f
C39 xb2_4.Y AVDD 0.541191f
C40 a_3612_3566# AVDD 0.35136f
C41 xa3.A VDD_ROSC 0.416232f
C42 xa3.Y a_2244_1806# 0.154165f
C43 xa3.A AVDD 0.952092f
C44 xb2_1.Y xb2_0.Y 0.196604f
C45 a_3612_3918# AVDD 0.35136f
C46 xa3.AN VDD_ROSC 0.413728f
C47 xb2_1.Y a_4764_2158# 0.126366f
C48 xa3.AN AVDD 0.828857f
C49 xb1.B VDD_ROSC 0.131663f
C50 xb1.B AVDD 0.635233f
C51 xa3.Y a_2244_2158# 0.140489f
C52 a_3612_4270# AVDD 0.35136f
C53 xb3.MP1.G AVDD 0.475974f
C54 xa3.YN xa3.xc2b.S 0.122641f
C55 a_3612_4622# AVDD 0.334453f
C56 xa3.AN a_1092_1102# 0.17278f
C57 xb2_2.Y xb2_1.Y 0.196604f
C58 xa3.YN xa3.Y 0.607411f
C59 xb2_2.Y a_4764_2510# 0.126366f
C60 AVDD PWRUP_1V8 0.751836f
C61 xa3.A a_1092_1806# 0.174769f
C62 xb1.B xb2_0.A 0.209066f
C63 AVDD CK 0.611632f
C64 AVDD VDD_ROSC 1.39916f
C65 a_3612_750# AVDD 0.335791f
C66 xb2_3.Y xb2_2.Y 0.196604f
C67 a_2244_750# AVDD 0.366882f
C68 xa3.A xa3.Y 0.293964f
C69 xb2_3.Y a_4764_2862# 0.126366f
C70 a_3612_1102# AVDD 0.352245f
C71 a_2244_1102# AVDD 0.363112f
C72 xa3.AN xa3.Y 0.192335f
C73 xa3.xc1b.S AVDD 0.152624f
C74 xa3.A xa3.YN 0.145399f
C75 a_3612_1454# AVDD 0.352245f
C76 PWRUP_1V8 AVSS 1.25525f
C77 CK AVSS 1.65304f
C78 VDD_ROSC AVSS 1.30035f
C79 AVDD AVSS 43.0788f
C80 a_4764_750# AVSS 0.492956f $ **FLOATING
C81 a_3612_750# AVSS 0.128212f $ **FLOATING
C82 a_2244_750# AVSS 0.127404f $ **FLOATING
C83 a_1092_750# AVSS 0.491389f $ **FLOATING
C84 a_4764_1102# AVSS 0.366247f $ **FLOATING
C85 a_1092_1102# AVSS 0.383754f $ **FLOATING
C86 xb1.MN1.S AVSS 0.175159f
C87 a_4764_1454# AVSS 0.380481f $ **FLOATING
C88 a_1092_1454# AVSS 0.388702f $ **FLOATING
C89 xb2_0.A AVSS 0.982003f
C90 a_4764_1806# AVSS 0.38397f $ **FLOATING
C91 a_1092_1806# AVSS 0.387701f $ **FLOATING
C92 xb2_0.Y AVSS 0.897154f
C93 a_4764_2158# AVSS 0.383938f $ **FLOATING
C94 a_1092_2158# AVSS 0.384097f $ **FLOATING
C95 xb2_1.Y AVSS 0.892951f
C96 xa3.Y AVSS 1.91185f
C97 xa4.Y AVSS 0.216345f
C98 a_4764_2510# AVSS 0.383925f $ **FLOATING
C99 a_1092_2510# AVSS 0.387855f $ **FLOATING
C100 xb2_2.Y AVSS 0.892866f
C101 xa3.YN AVSS 1.43322f
C102 a_4764_2862# AVSS 0.383917f $ **FLOATING
C103 a_1092_2862# AVSS 0.467284f $ **FLOATING
C104 xb2_3.Y AVSS 0.892823f
C105 a_4764_3214# AVSS 0.383831f $ **FLOATING
C106 a_1092_3214# AVSS 0.530885f $ **FLOATING
C107 xb2_4.Y AVSS 0.892662f
C108 a_4764_3566# AVSS 0.381065f $ **FLOATING
C109 xa3.A AVSS 3.21571f
C110 a_4764_3918# AVSS 0.381081f $ **FLOATING
C111 xa3.AN AVSS 3.84566f
C112 xb1.B AVSS 2.59951f
C113 a_4764_4270# AVSS 0.468519f $ **FLOATING
C114 xb3.MP1.G AVSS 0.118907f
C115 a_4764_4622# AVSS 0.567933f $ **FLOATING
C116 a_3612_4622# AVSS 0.128448f $ **FLOATING
.ends

